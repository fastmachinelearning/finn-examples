`timescale 1 ps / 1 ps

module TEMPLATE_design_wrapper
   (ddr3_sdram_addr,
    ddr3_sdram_ba,
    ddr3_sdram_cas_n,
    ddr3_sdram_ck_n,
    ddr3_sdram_ck_p,
    ddr3_sdram_cke,
    ddr3_sdram_cs_n,
    ddr3_sdram_dm,
    ddr3_sdram_dq,
    ddr3_sdram_dqs_n,
    ddr3_sdram_dqs_p,
    ddr3_sdram_odt,
    ddr3_sdram_ras_n,
    ddr3_sdram_reset_n,
    ddr3_sdram_we_n,
//    qspi_flash_io0_io,
//    qspi_flash_io1_io,
//    qspi_flash_io2_io,
//    qspi_flash_io3_io,
//    qspi_flash_sck_io,
//    qspi_flash_ss_io,
    reset,
    sys_clock,
    usb_uart_rxd,
    usb_uart_txd,
    usb_uart_rxd_debug,
    usb_uart_txd_debug    
    );
  output [13:0]ddr3_sdram_addr;
  output [2:0]ddr3_sdram_ba;
  output ddr3_sdram_cas_n;
  output [0:0]ddr3_sdram_ck_n;
  output [0:0]ddr3_sdram_ck_p;
  output [0:0]ddr3_sdram_cke;
  output [0:0]ddr3_sdram_cs_n;
  output [1:0]ddr3_sdram_dm;
  inout [15:0]ddr3_sdram_dq;
  inout [1:0]ddr3_sdram_dqs_n;
  inout [1:0]ddr3_sdram_dqs_p;
  output [0:0]ddr3_sdram_odt;
  output ddr3_sdram_ras_n;
  output ddr3_sdram_reset_n;
  output ddr3_sdram_we_n;
//  inout qspi_flash_io0_io;
//  inout qspi_flash_io1_io;
//  inout qspi_flash_io2_io;
//  inout qspi_flash_io3_io;
//  inout qspi_flash_sck_io;
//  inout qspi_flash_ss_io;
  input reset;
  input sys_clock;
  input usb_uart_rxd;
  output usb_uart_txd;
  output usb_uart_rxd_debug;
  output usb_uart_txd_debug;

  wire [13:0]ddr3_sdram_addr;
  wire [2:0]ddr3_sdram_ba;
  wire ddr3_sdram_cas_n;
  wire [0:0]ddr3_sdram_ck_n;
  wire [0:0]ddr3_sdram_ck_p;
  wire [0:0]ddr3_sdram_cke;
  wire [0:0]ddr3_sdram_cs_n;
  wire [1:0]ddr3_sdram_dm;
  wire [15:0]ddr3_sdram_dq;
  wire [1:0]ddr3_sdram_dqs_n;
  wire [1:0]ddr3_sdram_dqs_p;
  wire [0:0]ddr3_sdram_odt;
  wire ddr3_sdram_ras_n;
  wire ddr3_sdram_reset_n;
  wire ddr3_sdram_we_n;
//  wire qspi_flash_io0_i;
//  wire qspi_flash_io0_io;
//  wire qspi_flash_io0_o;
//  wire qspi_flash_io0_t;
//  wire qspi_flash_io1_i;
//  wire qspi_flash_io1_io;
//  wire qspi_flash_io1_o;
//  wire qspi_flash_io1_t;
//  wire qspi_flash_io2_i;
//  wire qspi_flash_io2_io;
//  wire qspi_flash_io2_o;
//  wire qspi_flash_io2_t;
//  wire qspi_flash_io3_i;
//  wire qspi_flash_io3_io;
//  wire qspi_flash_io3_o;
//  wire qspi_flash_io3_t;
//  wire qspi_flash_sck_i;
//  wire qspi_flash_sck_io;
//  wire qspi_flash_sck_o;
//  wire qspi_flash_sck_t;
//  wire qspi_flash_ss_i;
//  wire qspi_flash_ss_io;
//  wire qspi_flash_ss_o;
//  wire qspi_flash_ss_t;  
  wire reset;
  wire sys_clock;
  wire usb_uart_rxd;
  wire usb_uart_txd;
  wire usb_uart_rxd_debug;
  wire usb_uart_txd_debug;
  
  assign usb_uart_rxd_debug = usb_uart_rxd;
  assign usb_uart_txd = usb_uart_txd_debug;
  
  
//  IOBUF qspi_flash_io0_iobuf
//       (.I(qspi_flash_io0_o),
//        .IO(qspi_flash_io0_io),
//        .O(qspi_flash_io0_i),
//        .T(qspi_flash_io0_t));
//  IOBUF qspi_flash_io1_iobuf
//       (.I(qspi_flash_io1_o),
//        .IO(qspi_flash_io1_io),
//        .O(qspi_flash_io1_i),
//        .T(qspi_flash_io1_t));
//  IOBUF qspi_flash_io2_iobuf
//       (.I(qspi_flash_io2_o),
//        .IO(qspi_flash_io2_io),
//        .O(qspi_flash_io2_i),
//        .T(qspi_flash_io2_t));
//  IOBUF qspi_flash_io3_iobuf
//       (.I(qspi_flash_io3_o),
//        .IO(qspi_flash_io3_io),
//        .O(qspi_flash_io3_i),
//        .T(qspi_flash_io3_t));
//  IOBUF qspi_flash_sck_iobuf
//       (.I(qspi_flash_sck_o),
//        .IO(qspi_flash_sck_io),
//        .O(qspi_flash_sck_i),
//        .T(qspi_flash_sck_t));
//  IOBUF qspi_flash_ss_iobuf
//       (.I(qspi_flash_ss_o),
//        .IO(qspi_flash_ss_io),
//        .O(qspi_flash_ss_i),
//        .T(qspi_flash_ss_t));
  TEMPLATE_design TEMPLATE_design_i
       (.ddr3_sdram_addr(ddr3_sdram_addr),
        .ddr3_sdram_ba(ddr3_sdram_ba),
        .ddr3_sdram_cas_n(ddr3_sdram_cas_n),
        .ddr3_sdram_ck_n(ddr3_sdram_ck_n),
        .ddr3_sdram_ck_p(ddr3_sdram_ck_p),
        .ddr3_sdram_cke(ddr3_sdram_cke),
        .ddr3_sdram_cs_n(ddr3_sdram_cs_n),
        .ddr3_sdram_dm(ddr3_sdram_dm),
        .ddr3_sdram_dq(ddr3_sdram_dq),
        .ddr3_sdram_dqs_n(ddr3_sdram_dqs_n),
        .ddr3_sdram_dqs_p(ddr3_sdram_dqs_p),
        .ddr3_sdram_odt(ddr3_sdram_odt),
        .ddr3_sdram_ras_n(ddr3_sdram_ras_n),
        .ddr3_sdram_reset_n(ddr3_sdram_reset_n),
        .ddr3_sdram_we_n(ddr3_sdram_we_n),
//        .qspi_flash_io0_i(qspi_flash_io0_i),
//        .qspi_flash_io0_o(qspi_flash_io0_o),
//        .qspi_flash_io0_t(qspi_flash_io0_t),
//        .qspi_flash_io1_i(qspi_flash_io1_i),
//        .qspi_flash_io1_o(qspi_flash_io1_o),
//        .qspi_flash_io1_t(qspi_flash_io1_t),
//        .qspi_flash_io2_i(qspi_flash_io2_i),
//        .qspi_flash_io2_o(qspi_flash_io2_o),
//        .qspi_flash_io2_t(qspi_flash_io2_t),
//        .qspi_flash_io3_i(qspi_flash_io3_i),
//        .qspi_flash_io3_o(qspi_flash_io3_o),
//        .qspi_flash_io3_t(qspi_flash_io3_t),
//        .qspi_flash_sck_i(qspi_flash_sck_i),
//        .qspi_flash_sck_o(qspi_flash_sck_o),
//        .qspi_flash_sck_t(qspi_flash_sck_t),
//        .qspi_flash_ss_i(qspi_flash_ss_i),
//        .qspi_flash_ss_o(qspi_flash_ss_o),
//        .qspi_flash_ss_t(qspi_flash_ss_t),        
        .reset(reset),
        .sys_clock(sys_clock),
        .usb_uart_rxd(usb_uart_rxd),
        .usb_uart_txd_debug(usb_uart_txd_debug));
endmodule
